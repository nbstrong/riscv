-- A 32-bit RISC-V Processor
-- Nicholas Strong
--------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
--------------------------------------------------------------------------------
entity riscv is
    port (
        clkIn : in    std_logic;
        rstIn : in    std_logic
    );
end riscv;
--------------------------------------------------------------------------------
architecture behav of riscv is
    -- CONSTANTS ---------------------------------------------------------------
    -- SIGNALS -----------------------------------------------------------------
    -- ALIASES -----------------------------------------------------------------
    -- ATTRIBUTES --------------------------------------------------------------
begin
    -- PROGRAM COUNTER ---------------------------------------------------------
    p_counter_ent : entity work.prgcounter(behav)
        port map (
            clkIn       => clkIn,
            rstIn       => rstIn,
            addressOut  => address
        );

    -- PROGRAM MEM -------------------------------------------------------------
    -- REGISTERS ---------------------------------------------------------------
    -- ALU ---------------------------------------------------------------------
    -- DATA MEM ----------------------------------------------------------------
end behav;