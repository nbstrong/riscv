library IEEE;
use IEEE.std_logic_1164.all;
--------------------------------------------------------------------------------
entity register is
    port (
        clkIn : in    std_logic;
        rstIn : in    std_logic
    );
end register;
--------------------------------------------------------------------------------
architecture behav of register is
    -- CONSTANTS ---------------------------------------------------------------
    -- SIGNALS -----------------------------------------------------------------
    -- ALIASES -----------------------------------------------------------------
    -- ATTRIBUTES --------------------------------------------------------------
begin
    -- 32 registers of 64 bits
end behav;